module selector(inc_a, dec_a, inc_b, dec_b, inc_f, dec_f, sel, inc_pulse, dec_pulse, prev_pusle, next_pulse, clock);

output inc_a;
output dec_a;
output inc_b;
output dec_b;
output inc_f;
output dec_f;
output sel;

input inc_pulse;
input dec_pulse;
input prev_pusle;
input next_pulse;
input clock;

endmodule
